// Copyright (c) 2019 ETH Zurich, University of Bologna
//
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.

`ifndef AXI_TYPEDEF_SVH_
`define AXI_TYPEDEF_SVH_

`define AXI_TYPEDEF_AW_CHAN_T(aw_chan_t, addr_t, id_t, user_t)  \
  typedef struct packed {                                       \
    id_t              id;                                       \
    addr_t            addr;                                     \
    axi_pkg::len_t    len;                                      \
    axi_pkg::size_t   size;                                     \
    axi_pkg::burst_t  burst;                                    \
    logic             lock;                                     \
    axi_pkg::cache_t  cache;                                    \
    axi_pkg::prot_t   prot;                                     \
    axi_pkg::qos_t    qos;                                      \
    axi_pkg::region_t region;                                   \
    axi_pkg::atop_t   atop;                                     \
    user_t            user;                                     \
  } aw_chan_t;

`define AXI_TYPEDEF_W_CHAN_T(w_chan_t, data_t, strb_t, user_t)  \
  typedef struct packed {                                       \
    data_t data;                                                \
    strb_t strb;                                                \
    logic  last;                                                \
    user_t user;                                                \
  } w_chan_t;

`define AXI_TYPEDEF_B_CHAN_T(b_chan_t, id_t, user_t)  \
  typedef struct packed {                             \
    id_t            id;                               \
    axi_pkg::resp_t resp;                             \
    user_t          user;                             \
  } b_chan_t;

`define AXI_TYPEDEF_AR_CHAN_T(ar_chan_t, addr_t, id_t, user_t)  \
  typedef struct packed {                                       \
    id_t              id;                                       \
    addr_t            addr;                                     \
    axi_pkg::len_t    len;                                      \
    axi_pkg::size_t   size;                                     \
    axi_pkg::burst_t  burst;                                    \
    logic             lock;                                     \
    axi_pkg::cache_t  cache;                                    \
    axi_pkg::prot_t   prot;                                     \
    axi_pkg::qos_t    qos;                                      \
    axi_pkg::region_t region;                                   \
    user_t            user;                                     \
  } ar_chan_t;

`define AXI_TYPEDEF_R_CHAN_T(r_chan_t, data_t, id_t, user_t)  \
  typedef struct packed {                                     \
    id_t            id;                                       \
    data_t          data;                                     \
    axi_pkg::resp_t resp;                                     \
    logic           last;                                     \
    user_t          user;                                     \
  } r_chan_t;

`define AXI_TYPEDEF_REQ_T(req_t, aw_chan_t, w_chan_t, ar_chan_t)  \
  typedef struct packed {                                         \
    aw_chan_t aw;                                                 \
    logic     aw_valid;                                           \
    w_chan_t  w;                                                  \
    logic     w_valid;                                            \
    logic     b_ready;                                            \
    ar_chan_t ar;                                                 \
    logic     ar_valid;                                           \
    logic     r_ready;                                            \
  } req_t;

`define AXI_TYPEDEF_RESP_T(resp_t, b_chan_t, r_chan_t)  \
  typedef struct packed {                               \
    logic     aw_ready;                                 \
    logic     ar_ready;                                 \
    logic     w_ready;                                  \
    logic     b_valid;                                  \
    b_chan_t  b;                                        \
    logic     r_valid;                                  \
    r_chan_t  r;                                        \
  } resp_t;

// In AXI-Lite, the AR and AW channels have the same fields.
`define AXI_LITE_TYPEDEF_AX_CHAN_T(ax_chan_t, addr_t, id_t, user_t) \
  typedef struct packed {                                           \
    id_t              id;                                           \
    addr_t            addr;                                         \
    axi_pkg::size_t   size;                                         \
    axi_pkg::prot_t   prot;                                         \
    user_t            user;                                         \
  } ax_chan_t;

`define AXI_LITE_TYPEDEF_W_CHAN_T(w_chan_t, data_t, strb_t, user_t) \
  typedef struct packed {                                           \
    data_t data;                                                    \
    strb_t strb;                                                    \
    user_t user;                                                    \
  } w_chan_t;

`define AXI_LITE_TYPEDEF_B_CHAN_T(b_chan_t, id_t, user_t) \
  `AXI_TYPEDEF_B_CHAN_T(b_chan_t, id_t, user_t)

`define AXI_LITE_TYPEDEF_R_CHAN_T(r_chan_t, data_t, id_t, user_t) \
  typedef struct packed {                                         \
    id_t            id;                                           \
    data_t          data;                                         \
    axi_pkg::resp_t resp;                                         \
    user_t          user;                                         \
  } r_chan_t;

`define AXI_LITE_TYPEDEF_REQ_T(req_t, ax_chan_t, w_chan_t)  \
  typedef struct packed {                                   \
    ax_chan_t aw;                                           \
    logic     aw_valid;                                     \
    w_chan_t  w;                                            \
    logic     w_valid;                                      \
    logic     b_ready;                                      \
    ax_chan_t ar;                                           \
    logic     ar_valid;                                     \
    logic     r_ready;                                      \
  } req_t;

`define AXI_LITE_TYPEDEF_RESP_T(resp_t, b_chan_t, r_chan_t) \
  `AXI_TYPEDEF_RESP_T(resp_t, b_chan_t, r_chan_t)

`endif
