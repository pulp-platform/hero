// Copyright 2014-2018 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.

////////////////////////////////////////////////////////////////////////////////
// Company:        Institute of Integrated Systems // ETH Zurich              //
//                                                                            //
// Engineer:      Igor Loi - igor.loi@unibo.it                                //
//                                                                            //
// Additional contributions by:                                               //
//                 Davide Rossi                                               //
//                 Michael Gautschi                                           //
//                 Antonio Pullini                                            //
//                                                                            //
// Create Date:    12/03/2015                                                 //
// Design Name:    scm memory multiport                                       //
// Module Name:    register_file_2r_2w                                        //
// Project Name:   PULP                                                       //
// Language:       SystemVerilog                                              //
//                                                                            //
// Description:    scm memory multiport: 2 read Ports, 2 Write ports          //
//                                                                            //
// Revision:                                                                  //
// Revision v0.1 - File Created                                               //
// Revision v0.2 - Improved Identation                                        //
//                                                                            //
////////////////////////////////////////////////////////////////////////////////


module register_file_2r_2w_icache
#(
    parameter ADDR_WIDTH    = 5,
    parameter DATA_WIDTH    = 32
)
(
    // Clock and Reset
    input  logic                        clk,
    input  logic                        rst_n,

    input  logic                        test_en_i,

    //Read port R1
    input  logic                        ren_a_i,
    input  logic [ADDR_WIDTH-1:0]       raddr_a_i,
    output logic [DATA_WIDTH-1:0]       rdata_a_o,

    //Read port R2
    input  logic                        ren_b_i,
    input  logic [ADDR_WIDTH-1:0]       raddr_b_i,
    output logic [DATA_WIDTH-1:0]       rdata_b_o,

    // Write port W1
    input logic [ADDR_WIDTH-1:0]        waddr_a_i,
    input logic [DATA_WIDTH-1:0]        wdata_a_i,
    input logic                         we_a_i,

    // Write port W2
    input logic [ADDR_WIDTH-1:0]        waddr_b_i,
    input logic [DATA_WIDTH-1:0]        wdata_b_i,
    input logic                         we_b_i
);

    localparam    NUM_WORDS = 2**ADDR_WIDTH;

    // Read address register, located at the input of the address decoder
    logic [ADDR_WIDTH-1:0]                         RAddrRegxDPa;
    logic [ADDR_WIDTH-1:0]                         RAddrRegxDPb;
    logic [NUM_WORDS-1:0]                          RAddrOneHotxD;


    logic [DATA_WIDTH-1:0]                         MemContentxDP[NUM_WORDS];

    logic [NUM_WORDS-1:0]                          WAddrOneHotxDa;
    logic [NUM_WORDS-1:0]                          WAddrOneHotxDb;
    logic [NUM_WORDS-1:0]                          WAddrOneHotxDb_reg;

    logic [NUM_WORDS-1:0]                          ClocksxC;
`ifndef RF_2R2W_FF
    logic [DATA_WIDTH-1:0]                         WDataIntxDa;
    logic [DATA_WIDTH-1:0]                         WDataIntxDb;
`endif

    logic clk_int;

    logic we_int;

    int unsigned i;
    int unsigned j;
`ifndef RF_2R2W_FF
    int unsigned k;
`endif
    int unsigned l;
    int unsigned m;

    genvar x;
    genvar y;

    assign we_int = we_a_i | we_b_i;


    cluster_clock_gating CG_WE_GLOBAL
    (
        .clk_o(clk_int),
        .en_i(we_int),
        .test_en_i,
        .clk_i(clk)
    );

    //-----------------------------------------------------------------------------
    //-- READ : Read address register
    //-----------------------------------------------------------------------------

       always_ff @(posedge clk)
       begin : p_RAddrReg_a
               if(ren_a_i)
                       RAddrRegxDPa <= raddr_a_i;
       end

       always_ff @(posedge clk)
       begin : p_RAddrReg_b
               if(ren_b_i)
                       RAddrRegxDPb <= raddr_b_i;
       end

    //-----------------------------------------------------------------------------
    //-- READ : Read address decoder RAD
    //-----------------------------------------------------------------------------
    assign rdata_a_o = MemContentxDP[RAddrRegxDPa];
    assign rdata_b_o = MemContentxDP[RAddrRegxDPb];
    // assign rdata_a_o = MemContentxDP[raddr_a_i];
    // assign rdata_b_o = MemContentxDP[raddr_b_i];


    //-----------------------------------------------------------------------------
    //-- WRITE : Write Address Decoder (WAD), combinatorial process
    //-----------------------------------------------------------------------------
    always_comb
    begin : p_WADa
        for(i=0; i<NUM_WORDS; i++)
        begin : p_WordItera
            if ( (we_a_i == 1'b1 ) && (waddr_a_i == i) )
                    WAddrOneHotxDa[i] = 1'b1;
            else
                    WAddrOneHotxDa[i] = 1'b0;
        end
    end

    always_comb
    begin : p_WADb
        for(j=0; j<NUM_WORDS; j++)
        begin : p_WordIterb
            if ( (we_b_i == 1'b1 ) && (waddr_b_i == j) )
                    WAddrOneHotxDb[j] = 1'b1;
            else
                    WAddrOneHotxDb[j] = 1'b0;
        end
    end

    always_ff @(posedge clk_int)
    begin
        if(we_a_i | we_b_i)
            WAddrOneHotxDb_reg <= WAddrOneHotxDb;
    end

    //-----------------------------------------------------------------------------
    //-- WRITE : Clock gating (if integrated clock-gating cells are available)
    //-----------------------------------------------------------------------------
    generate
    for(x=0; x<NUM_WORDS; x++)
    begin : CG_CELL_WORD_ITER
        cluster_clock_gating CG_Inst
        (
            .clk_o(ClocksxC[x]),
            .en_i(WAddrOneHotxDa[x] | WAddrOneHotxDb[x]),
            .test_en_i,
            .clk_i(clk_int)
        );
    end
    endgenerate

`ifndef RF_2R2W_FF
    //-----------------------------------------------------------------------------
    // WRITE : SAMPLE INPUT DATA
    //---------------------------------------------------------------------------
    always_ff @(posedge clk)
    begin : sample_waddr
        if(we_a_i)
            WDataIntxDa <= wdata_a_i;
        if(we_b_i)
            WDataIntxDb <= wdata_b_i;
    end
`endif

    //-----------------------------------------------------------------------------
    //-- WRITE : Write operation
    //-----------------------------------------------------------------------------
    //-- Generate M = WORDS sequential processes, each of which describes one
    //-- word of the memory. The processes are synchronized with the clocks
    //-- ClocksxC(i), i = 0, 1, ..., M-1
    //-- Use active low, i.e. transparent on low latches as storage elements
    //-- Data is sampled on rising clock edge


`ifdef RF_2R2W_FF
    for (genvar k = 0; k < NUM_WORDS; k++) begin: gen_ff
      always_ff @(posedge ClocksxC[k]) begin
        if (WAddrOneHotxDb[k]) begin
          if (we_b_i) begin
            MemContentxDP[k] <= wdata_b_i;
          end
        `ifdef FPGA
        end
        if (WAddrOneHotxDa[k]) begin
        `else
        end else begin
        `endif
          if (we_a_i) begin
            MemContentxDP[k] <= wdata_a_i;
          end
        end
      end
    end
`else
    always_latch
    begin : latch_wdata
        for(k=0; k<NUM_WORDS; k++)
        begin : w_WordIter
            if( ClocksxC[k] == 1'b1)
                MemContentxDP[k] <= WAddrOneHotxDb_reg[k] ? WDataIntxDb : WDataIntxDa;
        end
    end
`endif

endmodule
